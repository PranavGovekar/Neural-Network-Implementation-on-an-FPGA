`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/27/2022 07:58:20 PM
// Design Name: 
// Module Name: neuron_256
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module neuron_256(input_weights_256,bias_256,out_256);

input signed [0:2047] input_weights_256;
input signed [7:0] bias_256;
output signed [31:0] out_256;

reg signed [8:0] image_array [0:255];
wire signed [7:0] weights_256 [0:255];

assign {weights_256[0],weights_256[1],weights_256[2],weights_256[3],weights_256[4],weights_256[5],weights_256[6],weights_256[7],weights_256[8],weights_256[9],weights_256[10],weights_256[11],weights_256[12],weights_256[13],weights_256[14],weights_256[15],weights_256[16],weights_256[17],weights_256[18],weights_256[19],weights_256[20],weights_256[21],weights_256[22],weights_256[23],weights_256[24],weights_256[25],weights_256[26],weights_256[27],weights_256[28],weights_256[29],weights_256[30],weights_256[31],weights_256[32],weights_256[33],weights_256[34],weights_256[35],weights_256[36],weights_256[37],weights_256[38],weights_256[39],weights_256[40],weights_256[41],weights_256[42],weights_256[43],weights_256[44],weights_256[45],weights_256[46],weights_256[47],weights_256[48],weights_256[49],weights_256[50],weights_256[51],weights_256[52],weights_256[53],weights_256[54],weights_256[55],weights_256[56],weights_256[57],weights_256[58],weights_256[59],weights_256[60],weights_256[61],weights_256[62],weights_256[63],weights_256[64],weights_256[65],weights_256[66],weights_256[67],weights_256[68],weights_256[69],weights_256[70],weights_256[71],weights_256[72],weights_256[73],weights_256[74],weights_256[75],weights_256[76],weights_256[77],weights_256[78],weights_256[79],weights_256[80],weights_256[81],weights_256[82],weights_256[83],weights_256[84],weights_256[85],weights_256[86],weights_256[87],weights_256[88],weights_256[89],weights_256[90],weights_256[91],weights_256[92],weights_256[93],weights_256[94],weights_256[95],weights_256[96],weights_256[97],weights_256[98],weights_256[99],weights_256[100],weights_256[101],weights_256[102],weights_256[103],weights_256[104],weights_256[105],weights_256[106],weights_256[107],weights_256[108],weights_256[109],weights_256[110],weights_256[111],weights_256[112],weights_256[113],weights_256[114],weights_256[115],weights_256[116],weights_256[117],weights_256[118],weights_256[119],weights_256[120],weights_256[121],weights_256[122],weights_256[123],weights_256[124],weights_256[125],weights_256[126],weights_256[127],weights_256[128],weights_256[129],weights_256[130],weights_256[131],weights_256[132],weights_256[133],weights_256[134],weights_256[135],weights_256[136],weights_256[137],weights_256[138],weights_256[139],weights_256[140],weights_256[141],weights_256[142],weights_256[143],weights_256[144],weights_256[145],weights_256[146],weights_256[147],weights_256[148],weights_256[149],weights_256[150],weights_256[151],weights_256[152],weights_256[153],weights_256[154],weights_256[155],weights_256[156],weights_256[157],weights_256[158],weights_256[159],weights_256[160],weights_256[161],weights_256[162],weights_256[163],weights_256[164],weights_256[165],weights_256[166],weights_256[167],weights_256[168],weights_256[169],weights_256[170],weights_256[171],weights_256[172],weights_256[173],weights_256[174],weights_256[175],weights_256[176],weights_256[177],weights_256[178],weights_256[179],weights_256[180],weights_256[181],weights_256[182],weights_256[183],weights_256[184],weights_256[185],weights_256[186],weights_256[187],weights_256[188],weights_256[189],weights_256[190],weights_256[191],weights_256[192],weights_256[193],weights_256[194],weights_256[195],weights_256[196],weights_256[197],weights_256[198],weights_256[199],weights_256[200],weights_256[201],weights_256[202],weights_256[203],weights_256[204],weights_256[205],weights_256[206],weights_256[207],weights_256[208],weights_256[209],weights_256[210],weights_256[211],weights_256[212],weights_256[213],weights_256[214],weights_256[215],weights_256[216],weights_256[217],weights_256[218],weights_256[219],weights_256[220],weights_256[221],weights_256[222],weights_256[223],weights_256[224],weights_256[225],weights_256[226],weights_256[227],weights_256[228],weights_256[229],weights_256[230],weights_256[231],weights_256[232],weights_256[233],weights_256[234],weights_256[235],weights_256[236],weights_256[237],weights_256[238],weights_256[239],weights_256[240],weights_256[241],weights_256[242],weights_256[243],weights_256[244],weights_256[245],weights_256[246],weights_256[247],weights_256[248],weights_256[249],weights_256[250],weights_256[251],weights_256[252],weights_256[253],weights_256[254],weights_256[255]} = input_weights_256;

initial
    begin
        $readmemb ("image0.mem", image_array);
    end
    
assign out_256 = ((image_array[0]*weights_256[0])+(image_array[1]*weights_256[1])+(image_array[2]*weights_256[2])+(image_array[3]*weights_256[3])+(image_array[4]*weights_256[4])+(image_array[5]*weights_256[5])+(image_array[6]*weights_256[6])+(image_array[7]*weights_256[7])+(image_array[8]*weights_256[8])+(image_array[9]*weights_256[9])+(image_array[10]*weights_256[10])+(image_array[11]*weights_256[11])+(image_array[12]*weights_256[12])+(image_array[13]*weights_256[13])+(image_array[14]*weights_256[14])+(image_array[15]*weights_256[15])+(image_array[16]*weights_256[16])+(image_array[17]*weights_256[17])+(image_array[18]*weights_256[18])+(image_array[19]*weights_256[19])+(image_array[20]*weights_256[20])+(image_array[21]*weights_256[21])+(image_array[22]*weights_256[22])+(image_array[23]*weights_256[23])+(image_array[24]*weights_256[24])+(image_array[25]*weights_256[25])+(image_array[26]*weights_256[26])+(image_array[27]*weights_256[27])+(image_array[28]*weights_256[28])+(image_array[29]*weights_256[29])+(image_array[30]*weights_256[30])+(image_array[31]*weights_256[31])+(image_array[32]*weights_256[32])+(image_array[33]*weights_256[33])+(image_array[34]*weights_256[34])+(image_array[35]*weights_256[35])+(image_array[36]*weights_256[36])+(image_array[37]*weights_256[37])+(image_array[38]*weights_256[38])+(image_array[39]*weights_256[39])+(image_array[40]*weights_256[40])+(image_array[41]*weights_256[41])+(image_array[42]*weights_256[42])+(image_array[43]*weights_256[43])+(image_array[44]*weights_256[44])+(image_array[45]*weights_256[45])+(image_array[46]*weights_256[46])+(image_array[47]*weights_256[47])+(image_array[48]*weights_256[48])+(image_array[49]*weights_256[49])+(image_array[50]*weights_256[50])+(image_array[51]*weights_256[51])+(image_array[52]*weights_256[52])+(image_array[53]*weights_256[53])+(image_array[54]*weights_256[54])+(image_array[55]*weights_256[55])+(image_array[56]*weights_256[56])+(image_array[57]*weights_256[57])+(image_array[58]*weights_256[58])+(image_array[59]*weights_256[59])+(image_array[60]*weights_256[60])+(image_array[61]*weights_256[61])+(image_array[62]*weights_256[62])+(image_array[63]*weights_256[63])+(image_array[64]*weights_256[64])+(image_array[65]*weights_256[65])+(image_array[66]*weights_256[66])+(image_array[67]*weights_256[67])+(image_array[68]*weights_256[68])+(image_array[69]*weights_256[69])+(image_array[70]*weights_256[70])+(image_array[71]*weights_256[71])+(image_array[72]*weights_256[72])+(image_array[73]*weights_256[73])+(image_array[74]*weights_256[74])+(image_array[75]*weights_256[75])+(image_array[76]*weights_256[76])+(image_array[77]*weights_256[77])+(image_array[78]*weights_256[78])+(image_array[79]*weights_256[79])+(image_array[80]*weights_256[80])+(image_array[81]*weights_256[81])+(image_array[82]*weights_256[82])+(image_array[83]*weights_256[83])+(image_array[84]*weights_256[84])+(image_array[85]*weights_256[85])+(image_array[86]*weights_256[86])+(image_array[87]*weights_256[87])+(image_array[88]*weights_256[88])+(image_array[89]*weights_256[89])+(image_array[90]*weights_256[90])+(image_array[91]*weights_256[91])+(image_array[92]*weights_256[92])+(image_array[93]*weights_256[93])+(image_array[94]*weights_256[94])+(image_array[95]*weights_256[95])+(image_array[96]*weights_256[96])+(image_array[97]*weights_256[97])+(image_array[98]*weights_256[98])+(image_array[99]*weights_256[99])+(image_array[100]*weights_256[100])+(image_array[101]*weights_256[101])+(image_array[102]*weights_256[102])+(image_array[103]*weights_256[103])+(image_array[104]*weights_256[104])+(image_array[105]*weights_256[105])+(image_array[106]*weights_256[106])+(image_array[107]*weights_256[107])+(image_array[108]*weights_256[108])+(image_array[109]*weights_256[109])+(image_array[110]*weights_256[110])+(image_array[111]*weights_256[111])+(image_array[112]*weights_256[112])+(image_array[113]*weights_256[113])+(image_array[114]*weights_256[114])+(image_array[115]*weights_256[115])+(image_array[116]*weights_256[116])+(image_array[117]*weights_256[117])+(image_array[118]*weights_256[118])+(image_array[119]*weights_256[119])+(image_array[120]*weights_256[120])+(image_array[121]*weights_256[121])+(image_array[122]*weights_256[122])+(image_array[123]*weights_256[123])+(image_array[124]*weights_256[124])+(image_array[125]*weights_256[125])+(image_array[126]*weights_256[126])+(image_array[127]*weights_256[127])+(image_array[128]*weights_256[128])+(image_array[129]*weights_256[129])+(image_array[130]*weights_256[130])+(image_array[131]*weights_256[131])+(image_array[132]*weights_256[132])+(image_array[133]*weights_256[133])+(image_array[134]*weights_256[134])+(image_array[135]*weights_256[135])+(image_array[136]*weights_256[136])+(image_array[137]*weights_256[137])+(image_array[138]*weights_256[138])+(image_array[139]*weights_256[139])+(image_array[140]*weights_256[140])+(image_array[141]*weights_256[141])+(image_array[142]*weights_256[142])+(image_array[143]*weights_256[143])+(image_array[144]*weights_256[144])+(image_array[145]*weights_256[145])+(image_array[146]*weights_256[146])+(image_array[147]*weights_256[147])+(image_array[148]*weights_256[148])+(image_array[149]*weights_256[149])+(image_array[150]*weights_256[150])+(image_array[151]*weights_256[151])+(image_array[152]*weights_256[152])+(image_array[153]*weights_256[153])+(image_array[154]*weights_256[154])+(image_array[155]*weights_256[155])+(image_array[156]*weights_256[156])+(image_array[157]*weights_256[157])+(image_array[158]*weights_256[158])+(image_array[159]*weights_256[159])+(image_array[160]*weights_256[160])+(image_array[161]*weights_256[161])+(image_array[162]*weights_256[162])+(image_array[163]*weights_256[163])+(image_array[164]*weights_256[164])+(image_array[165]*weights_256[165])+(image_array[166]*weights_256[166])+(image_array[167]*weights_256[167])+(image_array[168]*weights_256[168])+(image_array[169]*weights_256[169])+(image_array[170]*weights_256[170])+(image_array[171]*weights_256[171])+(image_array[172]*weights_256[172])+(image_array[173]*weights_256[173])+(image_array[174]*weights_256[174])+(image_array[175]*weights_256[175])+(image_array[176]*weights_256[176])+(image_array[177]*weights_256[177])+(image_array[178]*weights_256[178])+(image_array[179]*weights_256[179])+(image_array[180]*weights_256[180])+(image_array[181]*weights_256[181])+(image_array[182]*weights_256[182])+(image_array[183]*weights_256[183])+(image_array[184]*weights_256[184])+(image_array[185]*weights_256[185])+(image_array[186]*weights_256[186])+(image_array[187]*weights_256[187])+(image_array[188]*weights_256[188])+(image_array[189]*weights_256[189])+(image_array[190]*weights_256[190])+(image_array[191]*weights_256[191])+(image_array[192]*weights_256[192])+(image_array[193]*weights_256[193])+(image_array[194]*weights_256[194])+(image_array[195]*weights_256[195])+(image_array[196]*weights_256[196])+(image_array[197]*weights_256[197])+(image_array[198]*weights_256[198])+(image_array[199]*weights_256[199])+(image_array[200]*weights_256[200])+(image_array[201]*weights_256[201])+(image_array[202]*weights_256[202])+(image_array[203]*weights_256[203])+(image_array[204]*weights_256[204])+(image_array[205]*weights_256[205])+(image_array[206]*weights_256[206])+(image_array[207]*weights_256[207])+(image_array[208]*weights_256[208])+(image_array[209]*weights_256[209])+(image_array[210]*weights_256[210])+(image_array[211]*weights_256[211])+(image_array[212]*weights_256[212])+(image_array[213]*weights_256[213])+(image_array[214]*weights_256[214])+(image_array[215]*weights_256[215])+(image_array[216]*weights_256[216])+(image_array[217]*weights_256[217])+(image_array[218]*weights_256[218])+(image_array[219]*weights_256[219])+(image_array[220]*weights_256[220])+(image_array[221]*weights_256[221])+(image_array[222]*weights_256[222])+(image_array[223]*weights_256[223])+(image_array[224]*weights_256[224])+(image_array[225]*weights_256[225])+(image_array[226]*weights_256[226])+(image_array[227]*weights_256[227])+(image_array[228]*weights_256[228])+(image_array[229]*weights_256[229])+(image_array[230]*weights_256[230])+(image_array[231]*weights_256[231])+(image_array[232]*weights_256[232])+(image_array[233]*weights_256[233])+(image_array[234]*weights_256[234])+(image_array[235]*weights_256[235])+(image_array[236]*weights_256[236])+(image_array[237]*weights_256[237])+(image_array[238]*weights_256[238])+(image_array[239]*weights_256[239])+(image_array[240]*weights_256[240])+(image_array[241]*weights_256[241])+(image_array[242]*weights_256[242])+(image_array[243]*weights_256[243])+(image_array[244]*weights_256[244])+(image_array[245]*weights_256[245])+(image_array[246]*weights_256[246])+(image_array[247]*weights_256[247])+(image_array[248]*weights_256[248])+(image_array[249]*weights_256[249])+(image_array[250]*weights_256[250])+(image_array[251]*weights_256[251])+(image_array[252]*weights_256[252])+(image_array[253]*weights_256[253])+(image_array[254]*weights_256[254])+(image_array[255]*weights_256[255])+ bias_256);

endmodule
